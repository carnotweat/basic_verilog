module main;
  initial 
   begin
    $display("Learning Verilog is easy");
    $finish ;
   end
endmodule
